`define ALU_OP_MOVE 4'b0000 //move Rr to Rd
