
`define ALU_OP_COPY_TEST 	4'b0000
`define ALU_OP_COM 			4'b0001
`define ALU_OP_NEG 			4'b0010
`define ALU_OP_INC 			4'b0011
`define ALU_OP_DEC 			4'b0100
`define ALU_OP_SET_BIT 		4'b0101
`define ALU_OP_TRANSFERT 	4'b0111
`define ALU_OP_ADD 			4'b1001
`define ALU_OP_SUB 			4'b1010
`define ALU_OP_AND 			4'b1011
`define ALU_OP_OR 			4'b1100
`define ALU_OP_XOR 			4'b1101
`define ALU_OP_SWAP 		4'b1110
`define ALU_OP_RIGHT_SHIFT 	4'b1111

